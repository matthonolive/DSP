module fft #(parameter
  size = 1024
)(
  data_in,
  data_out
);



endmodule
